#include <stdio.h>



int main(void){
    char * mensaje = "Hola";


    printf("%s\n",mensaje);
    return 0;
    }
